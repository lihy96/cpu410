library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library work;
use work.constants.ALL;

entity fake_ram2 is
    Port ( 
           data_in, addr_in : in  STD_LOGIC_VECTOR (15 downto 0);
           --ram2OE, ram2WE, ram2EN: in std_logic;
		   RAM_READ_WRITE: in std_logic_vector(1 downto 0);
           data_out: out  STD_LOGIC_VECTOR (15 downto 0)
         );
end fake_ram2;

architecture Behavioral of fake_ram2 is
--type Inst_Array is array(11 downto 0) of std_logic_vector(15 downto 0);
--signal  ia: Inst_Array := 
signal ram2OE, ram2WE, ram2EN: std_logic;
begin
	ram2EN <= '0';
	ram2WE <= RAM_READ_WRITE(0);
	ram2OE <= not ram2WE;
	process(data_in, addr_in, ram_read_write)
	constant NOP: std_logic_vector(15 downto 0) := "0000100000000000";
	constant LI_R1_1: std_logic_vector(15 downto 0) := "0110100100000001";
	constant LI_R2_1: std_logic_vector(15 downto 0) := "0110101000000001";
	constant LI_R3_85: std_logic_vector(15 downto 0) := "0110101110000101";
	constant SLL_R3_R3_0: std_logic_vector(15 downto 0) := "0011001101100000";
	constant LI_R4_9: std_logic_vector(15 downto 0) := "0110110000001001";
	constant SW_R3_R1_0: std_logic_vector(15 downto 0) := "1101101100100000";
	constant SW_R3_R2_1: std_logic_vector(15 downto 0) := "1101101101000001";
	constant ADDU_R1_R2_R1: std_logic_vector(15 downto 0) := "1110000101000101";
	constant ADDU_R1_R2_R2: std_logic_vector(15 downto 0) := "1110000101001001";
	constant ADDIU_R3_2: std_logic_vector(15 downto 0) := "0100101100000010";
	constant ADDIU_R4_FF: std_logic_vector(15 downto 0) := "0100110011111111";
	constant BNEZ_R4_F9: std_logic_vector(15 downto 0) := "0010110011111001";
	begin
		if ram2OE = '0' and ram2EN = '0' then
			-- wait for 1 ns;
			case addr_in is
		when x"0000" =>
			data_out <= x"0000"; --ADDSP3 R0 0000
        when x"0001" =>
        	data_out <= x"0000"; --ADDSP3 R0 0000
        when x"0002" =>
        	data_out <= x"0800"; --NOP
        when x"0003" =>
        	data_out <= x"1061"; --B 0061
        when x"0004" =>
        	data_out <= x"0800"; --NOP
        when x"0005" =>
        	data_out <= x"0800"; --NOP
        when x"0006" =>
        	data_out <= x"0800"; --NOP
        when x"0007" =>
        	data_out <= x"0800"; --NOP
        when x"0008" =>
        	data_out <= x"6ebf"; --LI R6 00bf
        when x"0009" =>
        	data_out <= x"36c0"; --SLL R6 R6 0000
        when x"000a" =>
        	data_out <= x"4e10"; --ADDIU R6 0010
        when x"000b" =>
        	data_out <= x"de00"; --SW R6 R0 0000
        when x"000c" =>
        	data_out <= x"de21"; --SW R6 R1 0001
        when x"000d" =>
        	data_out <= x"de42"; --SW R6 R2 0002
        when x"000e" =>
        	data_out <= x"de84"; --SW R6 R4 0004
        when x"000f" =>
        	data_out <= x"dea5"; --SW R6 R5 0005
        when x"0010" =>
        	data_out <= x"9100"; --LW-SP R1 0000
        when x"0011" =>
        	data_out <= x"6301"; --ADDSP 0001
        when x"0012" =>
        	data_out <= x"68ff"; --LI R0 00ff
        when x"0013" =>
        	data_out <= x"e90c"; --AND R1 R0
        when x"0014" =>
        	data_out <= x"9200"; --LW-SP R2 0000
        when x"0015" =>
        	data_out <= x"6301"; --ADDSP 0001
        when x"0016" =>
        	data_out <= x"63ff"; --ADDSP ffff
        when x"0017" =>
        	data_out <= x"d300"; --SW-SP R3 0000
        when x"0018" =>
        	data_out <= x"63ff"; --ADDSP ffff
        when x"0019" =>
        	data_out <= x"d700"; --SW-SP R7 0000
        when x"001a" =>
        	data_out <= x"6b0f"; --LI R3 000f
        when x"001b" =>
        	data_out <= x"ef40"; --MFPC R7
        when x"001c" =>
        	data_out <= x"4f03"; --ADDIU R7 0003
        when x"001d" =>
        	data_out <= x"0800"; --NOP
        when x"001e" =>
        	data_out <= x"10ac"; --B 00ac
        when x"001f" =>
        	data_out <= x"0800"; --NOP
        when x"0020" =>
        	data_out <= x"6ebf"; --LI R6 00bf
        when x"0021" =>
        	data_out <= x"36c0"; --SLL R6 R6 0000
        when x"0022" =>
        	data_out <= x"de60"; --SW R6 R3 0000
        when x"0023" =>
        	data_out <= x"0800"; --NOP
        when x"0024" =>
        	data_out <= x"6ebf"; --LI R6 00bf
        when x"0025" =>
        	data_out <= x"36c0"; --SLL R6 R6 0000
        when x"0026" =>
        	data_out <= x"4e10"; --ADDIU R6 0010
        when x"0027" =>
        	data_out <= x"6800"; --LI R0 0000
        when x"0028" =>
        	data_out <= x"e82a"; --CMP R0 R1
        when x"0029" =>
        	data_out <= x"6102"; --BTNEZ 0002
        when x"002a" =>
        	data_out <= x"0800"; --NOP
        when x"002b" =>
        	data_out <= x"9e87"; --LW R6 R4 0007
        when x"002c" =>
        	data_out <= x"6820"; --LI R0 0020
        when x"002d" =>
        	data_out <= x"e82a"; --CMP R0 R1
        when x"002e" =>
        	data_out <= x"6102"; --BTNEZ 0002
        when x"002f" =>
        	data_out <= x"0800"; --NOP
        when x"0030" =>
        	data_out <= x"9e88"; --LW R6 R4 0008
        when x"0031" =>
        	data_out <= x"6810"; --LI R0 0010
        when x"0032" =>
        	data_out <= x"e82a"; --CMP R0 R1
        when x"0033" =>
        	data_out <= x"6102"; --BTNEZ 0002
        when x"0034" =>
        	data_out <= x"0800"; --NOP
        when x"0035" =>
        	data_out <= x"9e89"; --LW R6 R4 0009
        when x"0036" =>
        	data_out <= x"0800"; --NOP
        when x"0037" =>
        	data_out <= x"9ea6"; --LW R6 R5 0006
        when x"0038" =>
        	data_out <= x"eca2"; --SLT R4 R5
        when x"0039" =>
        	data_out <= x"610b"; --BTNEZ 000b
        when x"003a" =>
        	data_out <= x"0800"; --NOP
        when x"003b" =>
        	data_out <= x"de86"; --SW R6 R4 0006
        when x"003c" =>
        	data_out <= x"ef40"; --MFPC R7
        when x"003d" =>
        	data_out <= x"4f03"; --ADDIU R7 0003
        when x"003e" =>
        	data_out <= x"0800"; --NOP
        when x"003f" =>
        	data_out <= x"108b"; --B 008b
        when x"0040" =>
        	data_out <= x"0800"; --NOP
        when x"0041" =>
        	data_out <= x"6ebf"; --LI R6 00bf
        when x"0042" =>
        	data_out <= x"36c0"; --SLL R6 R6 0000
        when x"0043" =>
        	data_out <= x"de20"; --SW R6 R1 0000
        when x"0044" =>
        	data_out <= x"0800"; --NOP
        when x"0045" =>
        	data_out <= x"0800"; --NOP
        when x"0046" =>
        	data_out <= x"6b0f"; --LI R3 000f
        when x"0047" =>
        	data_out <= x"ef40"; --MFPC R7
        when x"0048" =>
        	data_out <= x"4f03"; --ADDIU R7 0003
        when x"0049" =>
        	data_out <= x"0800"; --NOP
        when x"004a" =>
        	data_out <= x"1080"; --B 0080
        when x"004b" =>
        	data_out <= x"0800"; --NOP
        when x"004c" =>
        	data_out <= x"6ebf"; --LI R6 00bf
        when x"004d" =>
        	data_out <= x"36c0"; --SLL R6 R6 0000
        when x"004e" =>
        	data_out <= x"de60"; --SW R6 R3 0000
        when x"004f" =>
        	data_out <= x"0800"; --NOP
        when x"0050" =>
        	data_out <= x"42c0"; --ADDIU3 R2 R6 0000
        when x"0051" =>
        	data_out <= x"f300"; --MFIH R3
        when x"0052" =>
        	data_out <= x"6880"; --LI R0 0080
        when x"0053" =>
        	data_out <= x"3000"; --SLL R0 R0 0000
        when x"0054" =>
        	data_out <= x"eb0d"; --OR R3 R0
        when x"0055" =>
        	data_out <= x"6fbf"; --LI R7 00bf
        when x"0056" =>
        	data_out <= x"37e0"; --SLL R7 R7 0000
        when x"0057" =>
        	data_out <= x"4f10"; --ADDIU R7 0010
        when x"0058" =>
        	data_out <= x"9f00"; --LW R7 R0 0000
        when x"0059" =>
        	data_out <= x"9f21"; --LW R7 R1 0001
        when x"005a" =>
        	data_out <= x"9f42"; --LW R7 R2 0002
        when x"005b" =>
        	data_out <= x"9f84"; --LW R7 R4 0004
        when x"005c" =>
        	data_out <= x"9fa5"; --LW R7 R5 0005
        when x"005d" =>
        	data_out <= x"9700"; --LW-SP R7 0000
        when x"005e" =>
        	data_out <= x"6301"; --ADDSP 0001
        when x"005f" =>
        	data_out <= x"6301"; --ADDSP 0001
        when x"0060" =>
        	data_out <= x"0800"; --NOP
        when x"0061" =>
        	data_out <= x"f301"; --MTIH R3
        when x"0062" =>
        	data_out <= x"ee00"; --JR R6
        when x"0063" =>
        	data_out <= x"93ff"; --LW-SP R3 00ff
        when x"0064" =>
        	data_out <= x"0800"; --NOP
        when x"0065" =>
        	data_out <= x"6807"; --LI R0 0007
        when x"0066" =>
        	data_out <= x"f001"; --MTIH R0
        when x"0067" =>
        	data_out <= x"68bf"; --LI R0 00bf
        when x"0068" =>
        	data_out <= x"3000"; --SLL R0 R0 0000
        when x"0069" =>
        	data_out <= x"4810"; --ADDIU R0 0010
        when x"006a" =>
        	data_out <= x"6400"; --MTSP R0
        when x"006b" =>
        	data_out <= x"0800"; --NOP
        when x"006c" =>
        	data_out <= x"6ebf"; --LI R6 00bf
        when x"006d" =>
        	data_out <= x"36c0"; --SLL R6 R6 0000
        when x"006e" =>
        	data_out <= x"4e10"; --ADDIU R6 0010
        when x"006f" =>
        	data_out <= x"6800"; --LI R0 0000
        when x"0070" =>
        	data_out <= x"de00"; --SW R6 R0 0000
        when x"0071" =>
        	data_out <= x"de01"; --SW R6 R0 0001
        when x"0072" =>
        	data_out <= x"de02"; --SW R6 R0 0002
        when x"0073" =>
        	data_out <= x"de03"; --SW R6 R0 0003
        when x"0074" =>
        	data_out <= x"de04"; --SW R6 R0 0004
        when x"0075" =>
        	data_out <= x"de05"; --SW R6 R0 0005
        when x"0076" =>
        	data_out <= x"de06"; --SW R6 R0 0006
        when x"0077" =>
        	data_out <= x"4801"; --ADDIU R0 0001
        when x"0078" =>
        	data_out <= x"de07"; --SW R6 R0 0007
        when x"0079" =>
        	data_out <= x"4801"; --ADDIU R0 0001
        when x"007a" =>
        	data_out <= x"de08"; --SW R6 R0 0008
        when x"007b" =>
        	data_out <= x"4801"; --ADDIU R0 0001
        when x"007c" =>
        	data_out <= x"de09"; --SW R6 R0 0009
        when x"007d" =>
        	data_out <= x"ef40"; --MFPC R7
        when x"007e" =>
        	data_out <= x"4f03"; --ADDIU R7 0003
        when x"007f" =>
        	data_out <= x"0800"; -- NOP
        when x"0080" =>
        	data_out <= x"104a"; -- B 004a
        when x"0081" =>
        	data_out <= x"6ebf"; -- LI R6 00bf
        when x"0082" =>
        	data_out <= x"36c0"; -- SLL R6 R6 0000
        when x"0083" =>
        	data_out <= x"684f"; -- LI R0 004f
        when x"0084" =>
        	data_out <= x"de00"; -- SW R6 R0 0000
        when x"0085" =>
        	data_out <= x"0800"; -- NOP
        when x"0086" =>
        	data_out <= x"ef40"; -- MFPC R7
        when x"0087" =>
        	data_out <= x"4f03"; -- ADDIU R7 0003
        when x"0088" =>
        	data_out <= x"0800"; -- NOP
        when x"0089" =>
        	data_out <= x"1041"; -- B 0041
        when x"008a" =>
        	data_out <= x"6ebf"; -- LI R6 00bf
        when x"008b" =>
        	data_out <= x"36c0"; -- SLL R6 R6 0000
        when x"008c" =>
        	data_out <= x"684b"; -- LI R0 004b
        when x"008d" =>
        	data_out <= x"de00"; -- SW R6 R0 0000
        when x"008e" =>
        	data_out <= x"0800"; -- NOP
        when x"008f" =>
        	data_out <= x"ef40"; -- MFPC R7
        when x"0090" =>
        	data_out <= x"4f03"; -- ADDIU R7 0003
        when x"0091" =>
        	data_out <= x"0800"; -- NOP
        when x"0092" =>
        	data_out <= x"1038"; -- B 0038
        when x"0093" =>
        	data_out <= x"6ebf"; -- LI R6 00bf
        when x"0094" =>
        	data_out <= x"36c0"; -- SLL R6 R6 0000
        when x"0095" =>
        	data_out <= x"680a"; -- LI R0 000a
        when x"0096" =>
        	data_out <= x"de00"; -- SW R6 R0 0000
        when x"0097" =>
        	data_out <= x"0800"; -- NOP
        when x"0098" =>
        	data_out <= x"ef40"; -- MFPC R7
        when x"0099" =>
        	data_out <= x"4f03"; -- ADDIU R7 0003
        when x"009a" =>
        	data_out <= x"0800"; -- NOP
        when x"009b" =>
        	data_out <= x"102f"; -- B 002f
        when x"009c" =>
        	data_out <= x"6ebf"; -- LI R6 00bf
        when x"009d" =>
        	data_out <= x"36c0"; -- SLL R6 R6 0000
        when x"009e" =>
        	data_out <= x"680d"; -- LI R0 000d
        when x"009f" =>
        	data_out <= x"de00"; -- SW R6 R0 0000
        when x"00a0" =>
        	data_out <= x"0800"; -- NOP
        when x"00a1" =>
        	data_out <= x"ef40"; -- MFPC R7
        when x"00a2" =>
        	data_out <= x"4f03"; -- ADDIU R7 0003
        when x"00a3" =>
        	data_out <= x"0800"; -- NOP
        when x"00a4" =>
        	data_out <= x"1031"; -- B 0031
        when x"00a5" =>
        	data_out <= x"0800"; -- NOP
        when x"00a6" =>
        	data_out <= x"6ebf"; -- LI R6 00bf
        when x"00a7" =>
        	data_out <= x"36c0"; -- SLL R6 R6 0000
        when x"00a8" =>
        	data_out <= x"9e20"; -- LW R6 R1 0000
        when x"00a9" =>
        	data_out <= x"6eff"; -- LI R6 00ff
        when x"00aa" =>
        	data_out <= x"e9cc"; -- AND R1 R6
        when x"00ab" =>
        	data_out <= x"0800"; -- NOP
        when x"00ac" =>
        	data_out <= x"6852"; -- LI R0 0052
        when x"00ad" =>
        	data_out <= x"e82a"; -- CMP R0 R1
        when x"00ae" =>
        	data_out <= x"6032"; -- BTEQZ 0032
        when x"00af" =>
        	data_out <= x"0800"; -- NOP
        when x"00b0" =>
        	data_out <= x"6844"; -- LI R0 0044
        when x"00b1" =>
        	data_out <= x"e82a"; -- CMP R0 R1
        when x"00b2" =>
        	data_out <= x"604d"; -- BTEQZ 004d
        when x"00b3" =>
        	data_out <= x"0800"; -- NOP
        when x"00b4" =>
        	data_out <= x"6841"; -- LI R0 0041
        when x"00b5" =>
        	data_out <= x"e82a"; -- CMP R0 R1
        when x"00b6" =>
        	data_out <= x"600e"; -- BTEQZ 000e
        when x"00b7" =>
        	data_out <= x"0800"; -- NOP
        when x"00b8" =>
        	data_out <= x"6855"; -- LI R0 0055
        when x"00b9" =>
        	data_out <= x"e82a"; -- CMP R0 R1
        when x"00ba" =>
        	data_out <= x"6007"; -- BTEQZ 0007
        when x"00bb" =>
        	data_out <= x"0800"; -- NOP
        when x"00bc" =>
        	data_out <= x"6847"; -- LI R0 0047
        when x"00bd" =>
        	data_out <= x"e82a"; -- CMP R0 R1
        when x"00be" =>
        	data_out <= x"6009"; -- BTEQZ 0009
        when x"00bf" =>
        	data_out <= x"0800"; -- NOP
        when x"00c0" =>
        	data_out <= x"17e0"; -- B ffe0
        when x"00c1" =>
        	data_out <= x"0800"; -- NOP
        when x"00c2" =>
        	data_out <= x"0800"; -- NOP
        when x"00c3" =>
        	data_out <= x"10c0"; -- B 00c0
        when x"00c4" =>
        	data_out <= x"0800"; -- NOP
        when x"00c5" =>
        	data_out <= x"0800"; -- NOP
        when x"00c6" =>
        	data_out <= x"1082"; -- B 0082
        when x"00c7" =>
        	data_out <= x"0800"; -- NOP
        when x"00c8" =>
        	data_out <= x"0800"; -- NOP
        when x"00c9" =>
        	data_out <= x"1103"; -- B 0103
        when x"00ca" =>
        	data_out <= x"0800"; -- NOP
        when x"00cb" =>
        	data_out <= x"0800"; -- NOP
        when x"00cc" =>
        	data_out <= x"6ebf"; -- LI R6 00bf
        when x"00cd" =>
        	data_out <= x"36c0"; -- SLL R6 R6 0000
        when x"00ce" =>
        	data_out <= x"4e01"; -- ADDIU R6 0001
        when x"00cf" =>
        	data_out <= x"9e00"; -- LW R6 R0 0000
        when x"00d0" =>
        	data_out <= x"6e01"; -- LI R6 0001
        when x"00d1" =>
        	data_out <= x"e8cc"; -- AND R0 R6
        when x"00d2" =>
        	data_out <= x"20f8"; -- BEQZ R0 fff8
        when x"00d3" =>
        	data_out <= x"0800"; -- NOP
        when x"00d4" =>
        	data_out <= x"ef00"; -- JR R7
        when x"00d5" =>
        	data_out <= x"0800"; -- NOP
        when x"00d6" =>
        	data_out <= x"0800"; -- NOP
        when x"00d7" =>
        	data_out <= x"6ebf"; -- LI R6 00bf
        when x"00d8" =>
        	data_out <= x"36c0"; -- SLL R6 R6 0000
        when x"00d9" =>
        	data_out <= x"4e01"; -- ADDIU R6 0001
        when x"00da" =>
        	data_out <= x"9e00"; -- LW R6 R0 0000
        when x"00db" =>
        	data_out <= x"6e02"; -- LI R6 0002
        when x"00dc" =>
        	data_out <= x"e8cc"; -- AND R0 R6
        when x"00dd" =>
        	data_out <= x"20f8"; -- BEQZ R0 fff8
        when x"00de" =>
        	data_out <= x"0800"; -- NOP
        when x"00df" =>
        	data_out <= x"ef00"; -- JR R7
        when x"00e0" =>
        	data_out <= x"0800"; -- NOP
        when x"00e1" =>
        	data_out <= x"6906"; -- LI R1 0006
        when x"00e2" =>
        	data_out <= x"6a06"; -- LI R2 0006
        when x"00e3" =>
        	data_out <= x"68bf"; -- LI R0 00bf
        when x"00e4" =>
        	data_out <= x"3000"; -- SLL R0 R0 0000
        when x"00e5" =>
        	data_out <= x"4810"; -- ADDIU R0 0010
        when x"00e6" =>
        	data_out <= x"e22f"; -- SUBU R2 R1 R3
        when x"00e7" =>
        	data_out <= x"e061"; -- ADDU R0 R3 R0
        when x"00e8" =>
        	data_out <= x"9860"; -- LW R0 R3 0000
        when x"00e9" =>
        	data_out <= x"ef40"; -- MFPC R7
        when x"00ea" =>
        	data_out <= x"4f03"; -- ADDIU R7 0003
        when x"00eb" =>
        	data_out <= x"0800"; -- NOP
        when x"00ec" =>
        	data_out <= x"17de"; -- B ffde
        when x"00ed" =>
        	data_out <= x"0800"; -- NOP
        when x"00ee" =>
        	data_out <= x"6ebf"; -- LI R6 00bf
        when x"00ef" =>
        	data_out <= x"36c0"; -- SLL R6 R6 0000
        when x"00f0" =>
        	data_out <= x"de60"; -- SW R6 R3 0000
        when x"00f1" =>
        	data_out <= x"3363"; -- SRA R3 R3 0000
        when x"00f2" =>
        	data_out <= x"ef40"; -- MFPC R7
        when x"00f3" =>
        	data_out <= x"4f03"; -- ADDIU R7 0003
        when x"00f4" =>
        	data_out <= x"0800"; -- NOP
        when x"00f5" =>
        	data_out <= x"17d5"; -- B ffd5
        when x"00f6" =>
        	data_out <= x"0800"; -- NOP
        when x"00f7" =>
        	data_out <= x"6ebf"; -- LI R6 00bf
        when x"00f8" =>
        	data_out <= x"36c0"; -- SLL R6 R6 0000
        when x"00f9" =>
        	data_out <= x"de60"; -- SW R6 R3 0000
        when x"00fa" =>
        	data_out <= x"49ff"; -- ADDIU R1 ffff
        when x"00fb" =>
        	data_out <= x"0800"; -- NOP
        when x"00fc" =>
        	data_out <= x"29e6"; -- BNEZ R1 ffe6
        when x"00fd" =>
        	data_out <= x"0800"; -- NOP
        when x"00fe" =>
        	data_out <= x"17a2"; -- B ffa2
        when x"00ff" =>
        	data_out <= x"0800"; -- NOP
        when x"0100" =>
        	data_out <= x"ef40"; -- MFPC R7
        when x"0101" =>
        	data_out <= x"4f03"; -- ADDIU R7 0003
        when x"0102" =>
        	data_out <= x"0800"; -- NOP
        when x"0103" =>
        	data_out <= x"17d2"; -- B ffd2
        when x"0104" =>
        	data_out <= x"0800"; -- NOP
        when x"0105" =>
        	data_out <= x"6ebf"; -- LI R6 00bf
        when x"0106" =>
        	data_out <= x"36c0"; -- SLL R6 R6 0000
        when x"0107" =>
        	data_out <= x"9ea0"; -- LW R6 R5 0000
        when x"0108" =>
        	data_out <= x"6eff"; -- LI R6 00ff
        when x"0109" =>
        	data_out <= x"edcc"; -- AND R5 R6
        when x"010a" =>
        	data_out <= x"0800"; -- NOP
        when x"010b" =>
        	data_out <= x"ef40"; -- MFPC R7
        when x"010c" =>
        	data_out <= x"4f03"; -- ADDIU R7 0003
        when x"010d" =>
        	data_out <= x"0800"; -- NOP
        when x"010e" =>
        	data_out <= x"17c7"; -- B ffc7
        when x"010f" =>
        	data_out <= x"0800"; -- NOP
        when x"0110" =>
        	data_out <= x"6ebf"; -- LI R6 00bf
        when x"0111" =>
        	data_out <= x"36c0"; -- SLL R6 R6 0000
        when x"0112" =>
        	data_out <= x"9e20"; -- LW R6 R1 0000
        when x"0113" =>
        	data_out <= x"6eff"; -- LI R6 00ff
        when x"0114" =>
        	data_out <= x"e9cc"; -- AND R1 R6
        when x"0115" =>
        	data_out <= x"0800"; -- NOP
        when x"0116" =>
        	data_out <= x"3120"; -- SLL R1 R1 0000
        when x"0117" =>
        	data_out <= x"e9ad"; -- OR R1 R5
        when x"0118" =>
        	data_out <= x"ef40"; -- MFPC R7
        when x"0119" =>
        	data_out <= x"4f03"; -- ADDIU R7 0003
        when x"011a" =>
        	data_out <= x"0800"; -- NOP
        when x"011b" =>
        	data_out <= x"17ba"; -- B ffba
        when x"011c" =>
        	data_out <= x"0800"; -- NOP
        when x"011d" =>
        	data_out <= x"6ebf"; -- LI R6 00bf
        when x"011e" =>
        	data_out <= x"36c0"; -- SLL R6 R6 0000
        when x"011f" =>
        	data_out <= x"9ea0"; -- LW R6 R5 0000
				--when "0000000000000000" =>
				--	data_out <= NOP;
				--when x"0001" => 
				    --data_out <= x"6c48";-- LI R4 0048
				--when x"0002" => 
				--    data_out <= x"6d85";-- LI R5 0085
				--when x"0003" => 
				--    data_out <= x"35a0";-- SLL R5 R5 0000
				--when x"0004" => 
				--    data_out <= x"6800";-- LI R0 0000
				--when x"0005" => 
				--    data_out <= x"6901";-- LI R1 0001
				--when x"0006" => 
				--    data_out <= x"dd00";-- SW R5 R0 0000
				--when x"0007" => 
				--    data_out <= x"dd01";-- SW R5 R0 0001
				--when x"0008" => 
				--    data_out <= x"dd22";-- SW R5 R1 0002
				--when x"0009" => 
				--    data_out <= x"4d03";-- ADDIU R5 0003
				--when x"000a" => 
				--    data_out <= x"dd00";-- SW R5 R0 0000
				--when x"000b" => 
				--    data_out <= x"dd01";-- SW R5 R0 0001
				--when x"000c" => 
				--    data_out <= x"dd22";-- SW R5 R1 0002
				--when x"000d" => 
				--    data_out <= x"4d03";-- ADDIU R5 0003
				--when x"000e" => 
				--    data_out <= x"9d1f";-- LW R5 R0 ffff
				--when x"000f" => 
				--    data_out <= x"9d3c";-- LW R5 R1 fffc
				--when x"0010" => 
				--    data_out <= x"e029";-- ADDU R0 R1 R2
				--when x"0011" => 
				--    data_out <= x"dd42";-- SW R5 R2 0002
				--when x"0012" => 
				--    data_out <= x"ea03";-- SLTU R2 R0
				--when x"0013" => 
				--    data_out <= x"6107";-- BTNEZ 0007
				--when x"0014" => 
				--    data_out <= x"0800";-- NOP
				--when x"0015" => 
				--    data_out <= x"ea23";-- SLTU R2 R1
				--when x"0016" => 
				--    data_out <= x"6104";-- BTNEZ 0004
				--when x"0017" => 
				--    data_out <= x"0800";-- NOP
				--when x"0018" => 
				--    data_out <= x"6b00";-- LI R3 0000
				--when x"0019" => 
				--    data_out <= x"1002";-- B 0002
				--when x"001a" => 
				--    data_out <= x"0800";-- NOP
				--when x"001b" => 
				--    data_out <= x"6b01";-- LI R3 0001
				--when x"001c" => 
				--    data_out <= x"9d1e";-- LW R5 R0 fffe
				--when x"001d" => 
				--    data_out <= x"9d3b";-- LW R5 R1 fffb
				--when x"001e" => 
				--    data_out <= x"e029";-- ADDU R0 R1 R2
				--when x"001f" => 
				--    data_out <= x"e349";-- ADDU R3 R2 R2
				--when x"0020" => 
				--    data_out <= x"dd41";-- SW R5 R2 0001
				--when x"0021" => 
				--    data_out <= x"ea03";-- SLTU R2 R0
				--when x"0022" => 
				--    data_out <= x"6107";-- BTNEZ 0007
				--when x"0023" => 
				--    data_out <= x"0800";-- NOP
				--when x"0024" => 
				--    data_out <= x"ea23";-- SLTU R2 R1
				--when x"0025" => 
				--    data_out <= x"6104";-- BTNEZ 0004
				--when x"0026" => 
				--    data_out <= x"0800";-- NOP
				--when x"0027" => 
				--    data_out <= x"6b00";-- LI R3 0000
				--when x"0028" => 
				--    data_out <= x"1002";-- B 0002
				--when x"0029" => 
				--    data_out <= x"0800";-- NOP
				--when x"002a" => 
				--    data_out <= x"6b01";-- LI R3 0001
				--when x"002b" => 
				--    data_out <= x"9d1d";-- LW R5 R0 fffd
				--when x"002c" => 
				--    data_out <= x"9d3a";-- LW R5 R1 fffa
				--when x"002d" => 
				--    data_out <= x"e029";-- ADDU R0 R1 R2
				--when x"002e" => 
				--    data_out <= x"e349";-- ADDU R3 R2 R2
				--when x"002f" => 
				--    data_out <= x"dd40";-- SW R5 R2 0000
				--when x"0030" => 
				--    data_out <= x"4cff";-- ADDIU R4 ffff
				--when x"0031" => 
				--    data_out <= x"4d03";-- ADDIU R5 0003
				--when x"0032" => 
				--    data_out <= x"2cdb";-- BNEZ R4 ffdb
				--when x"0033" => 
				--    data_out <= x"0800";-- NOP
				--when x"0034" => 
				--    data_out <= x"ffff";-- RET
				--when x"0035" => 
				--    data_out <= x"0800";-- NOP
				--when "0000000000000001" => 
				--	data_out <= LI_R1_1;
				--when "0000000000000010" => 
				--	data_out <= LI_R2_1;
				--when "0000000000000011" => 
				--	data_out <= LI_R3_85;
				--when "0000000000000100" => 
				--	data_out <= SLL_R3_R3_0;
				--when "0000000000000101" => 
				--	data_out <= LI_R4_9;
				--when "0000000000000110" => 
				--	data_out <= SW_R3_R1_0;
				--when "0000000000000111" => 
				--	data_out <= SW_R3_R2_1;
				--when "0000000000001000" => 
				--	data_out <= ADDU_R1_R2_R1;
				--when "0000000000001001" => 
				--	data_out <= ADDU_R1_R2_R2;
				--when "0000000000001010" => 
				--	data_out <= ADDIU_R3_2;
				--when "0000000000001011" => 
				--	data_out <= ADDIU_R4_FF;
				--when "0000000000001100" => 
				--	data_out <= BNEZ_R4_F9;
				--when "0000000000001101" =>
				--	data_out <= NOP;

				when others =>
					data_out <= NOP;
			end case ;
		end if;
	end process ;
end Behavioral;
