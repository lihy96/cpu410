library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.constants.all;

entity forward is
  port (
  	reg_bus: in std_logic_vector(11 downto 0) ;
 	reg_prev1: in std_logic_vector(3 downto 0) ;
 	reg_prev2: in std_logic_vector(3 downto 0) ;
 	
  ) ;
end entity ; -- forward

architecture Behavioral of forward is
	signal 

begin

end architecture ; -- Behavioral